LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY indexed_data IS
	PORT(
		op_code : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		res : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
	);
END ENTITY;

ARCHITECTURE bhr OF indexed_data IS
BEGIN
	PROCESS(op_code)
	BEGIN
	
	END PROCESS;
END ARCHITECTURE;
