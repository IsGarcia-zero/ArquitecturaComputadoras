library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
entity comparador16 is
    port (
        x, y: in std_logic_vector(15 downto 0);
        g0, l0: in std_logic;
        gtt, eqq, ltt: out std_logic
    );
end entity comparador16;

architecture Behavioral of comparador16 is
    signal gts, eqs, lts: std_logic_vector(1 downto 0);
    component comparador8 is
        port (
            x, y: in std_logic_vector(7 downto 0);
				g0, l0: in std_logic;
				gtt, eqq, ltt: out std_logic
        );
    end component comparador8;
begin
    comp0: comparador8 port map(x(7 downto 0), y(7 downto 0), g0, l0, gts(0), lts(0), eqs(0));
    comp1: comparador8 port map(x(15 downto 8), y(15 downto 8), gts(0), lts(0), gtt, eqq, ltt);
end architecture Behavioral;