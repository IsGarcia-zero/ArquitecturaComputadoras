LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC.UNSIGNED.ALL;

ENTITY stack IS
	PORT(
		input : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		clk : IN STD_LOGIC;
		push, pop; IN STD_LOGIC;
		sal : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE bhr OF stack IS
	SIGNAL i : INTEGER RANGE 0 TO 99 := 0;
	TYPE data IS ARRAY(99 DOWNTO 0) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL ram IS data;
BEGIN
	PROCESS(clk)
	BEGIN
		IF (RISING_EDGE(clk)) THEN
			IF(push = '1') THEN
				data(i) <= input;
				i <= i + 1;
			END ENTITY;
			IF(pop = '1' AND i > 0) THEN
				data(i) <= "0000000000000000";
				i <= i - 1;
			END ENTITY
		END ENTITY
	END PROCESS;
	



END ARCHITECTURE;