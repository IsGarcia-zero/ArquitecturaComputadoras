LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY join IS
	PORT(
		a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		b : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		enable : IN STD_LOGIC;
		ins : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		sal : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE bhr OF join IS
BEGIN
	WITH enable SELECT sal <=
		ins WHEN '1',
		b & a(11 DOWNTO 0) WHEN '0';
END ARCHITECTURE;

